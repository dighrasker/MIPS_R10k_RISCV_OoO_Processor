module ROB (
    input ROB_ENTRY_PACKET rob_entry;

    input   


    output RETIREMENT_PACKET retire_packet;
)