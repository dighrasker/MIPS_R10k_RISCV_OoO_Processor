`include "verilog/sys_defs.svh"

module 