`include "sys_defs.svh"

module Issue # (
) (
    // ------------- FROM FREDDY -------------- //
    input logic  [`PHYS_REG_SZ_R10K-1:0] complete_list_copy,

);

endmodule